
//design code goes here

module dut();



endmodule;
